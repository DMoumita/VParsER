module M;

time  b[2:0]=2;

endmodule
