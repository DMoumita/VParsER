module M;

reg [1:0] a, b = 1;

endmodule
