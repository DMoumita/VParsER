module M;

realtime  b[2:0]=2;

endmodule
