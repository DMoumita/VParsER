module m;

wand  w1;
wand  signed w7;
wand  w11[2:0];
wand  signed w9[2:0];
wand  wm21,w211[3:0],w4;
wand  w281[4:0],w21[9:3];

wand  signed n1,n2[3:0],n3;
wand  vectored [4:0] n5[2:0];
wand  scalared signed [4:0] nw9[2:0];
endmodule
