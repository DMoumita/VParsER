module M;

endmodule
