module M();
endmodule
