module M;

integer  a,b;
integer  x=1,y=2;
integer  x1[1:0],y1[2:1];
integer  xx1[1:0],yy1, z1[3:0],p=2;
endmodule
