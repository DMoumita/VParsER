module M;

realtime  a,b;
realtime  x=1,y=2;
realtime  x1[1:0],y1[2:1];
realtime  xx1[1:0],yy1, z1[3:0],p=2;
endmodule
