module M;

real  b[2:0]=2;

endmodule
