module M(input a, output b, input c);
endmodule
