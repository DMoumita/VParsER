module M(a);
input a;
endmodule
