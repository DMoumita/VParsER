module m;

trior  w1;
trior  signed w7;
trior  w11[2:0];
trior  signed w9[2:0];
trior  wm21,w211[3:0],w4;
trior  w281[4:0],w21[9:3];

trior  signed n1,n2[3:0],n3;
trior  vectored [4:0] n5[2:0];
trior  scalared signed [4:0] nw9[2:0];
endmodule
