module M;
  wire w1 = 1'b1;
  assign w2 = w1;
endmodule
