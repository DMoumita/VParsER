module M;

realtime [2:0 b;

endmodule
