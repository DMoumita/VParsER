module m;

tri1  w1;
tri1  signed w7;
tri1  w11[2:0];
tri1  signed w9[2:0];
tri1  wm21,w211[3:0],w4;
tri1  w281[4:0],w21[9:3];

tri1  signed n1,n2[3:0],n3;
tri1  vectored [4:0] n5[2:0];
tri1  scalared signed [4:0] nw9[2:0];
endmodule
