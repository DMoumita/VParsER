module M;
  wire w1 = 1'b1;
endmodule
