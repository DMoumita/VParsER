module M;

reg [1:0] b[2:0]=1;

endmodule
