module m;

tri0  w1;
tri0  signed w7;
tri0  w11[2:0];
tri0  signed w9[2:0];
tri0  wm21,w211[3:0],w4;
tri0  w281[4:0],w21[9:3];

tri0  signed n1,n2[3:0],n3;
tri0  vectored [4:0] n5[2:0];
tri0  scalared signed [4:0] nw9[2:0];
endmodule
