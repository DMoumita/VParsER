module M;

real [1:0] b[2:0]=2;

endmodule
