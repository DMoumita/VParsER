module M;
  wire (strong1, pull0) w1 = 1'b1;
endmodule
