module m;

wire    n5[2:0] =1'b0;
endmodule
