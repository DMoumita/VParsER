module m;

wire  w1;
wire  signed w7;
wire  w11[2:0];
wire  signed w9[2:0];
wire  wm21,w211[3:0],w4;
wire  w281[4:0],w21[9:3];

wire  signed n1,n2[3:0],n3;
wire  vectored [4:0] n5[2:0];
wire  scalared signed [4:0] nw9[2:0];
wire [4:0] m1;
wire [4:0] m2[2:0];
wire [4:0] m3[2:0],m4;
wire [4:0] m5[2:0],m41[5:1];
endmodule
