module m;

wor  w1;
wor  signed w7;
wor  w11[2:0];
wor  signed w9[2:0];
wor  wm21,w211[3:0],w4;
wor  w281[4:0],w21[9:3];

wor  signed n1,n2[3:0],n3;
wor  vectored [4:0] n5[2:0];
wor  scalared signed [4:0] nw9[2:0];
endmodule
