module m;

tri  w1;
tri  signed w7;
tri  w11[2:0];
tri  signed w9[2:0];
tri  wm21,w211[3:0],w4;
tri  w281[4:0],w21[9:3];

tri  signed n1,n2[3:0],n3;
tri  vectored [4:0] n5[2:0];
tri  scalared signed [4:0] nw9[2:0];
endmodule
