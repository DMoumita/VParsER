module M;

integer [2:0 b;

endmodule
