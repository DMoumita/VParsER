module M;

integer  b[2:0]=2;

endmodule
