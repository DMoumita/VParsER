module M;

time  a,b;
time  x=1,y=2;
time  x1[1:0],y1[2:1];
time  xx1[1:0],yy1, z1[3:0],p=2;
endmodule
