module M;

real [2:0 b;

endmodule
