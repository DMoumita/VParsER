module M(a);
endmodule
