module M(a,b,c);
input a;
output reg b;
wire a;
output time c;
endmodule
