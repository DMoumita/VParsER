module m;

wire   vectored n5[2:0];
endmodule
