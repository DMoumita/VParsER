module M;

real  a,b;
real  x=1,y=2;
real  x1[1:0],y1[2:1];
real  xx1[1:0],yy1, z1[3:0],p=2;
endmodule
