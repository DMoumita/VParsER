module m;

supply0  w1;
supply1  signed w7;
supply0  w11[2:0];
supply0  signed w9[2:0];
supply1  wm21,w211[3:0],w4;
supply1  w281[4:0],w21[9:3];

supply0  signed n1,n2[3:0],n3;
supply0  vectored [4:0] n5[2:0];
supply1  scalared signed [4:0] nw9[2:0];
supply1 [4:0] m1;
supply1 [4:0] m2[2:0];
supply1 [4:0] m3[2:0],m4;
supply0 [4:0] m5[2:0],m41[5:1];
endmodule
