module M;

time [1:0] b[2:0]=2;

endmodule
