module M;

time [2:0 b;

endmodule
