module M;

reg b[1:0][2:0]=1;

endmodule
