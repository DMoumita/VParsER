module m;

uwire  w1;
uwire  signed w7;
uwire  w11[2:0];
uwire  signed w9[2:0];
uwire  wm21,w211[3:0],w4;
uwire  w281[4:0],w21[9:3];

uwire  signed n1,n2[3:0],n3;
uwire  vectored [4:0] n5[2:0];
uwire  scalared signed [4:0] nw9[2:0];
endmodule
