module m;

wire (strong1, pull0) w1;

endmodule
