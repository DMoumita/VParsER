module m;

triand  w1;
triand  signed w7;
triand  w11[2:0];
triand  signed w9[2:0];
triand  wm21,w211[3:0],w4;
triand  w281[4:0],w21[9:3];

triand  signed n1,n2[3:0],n3;
triand  vectored [4:0] n5[2:0];
triand  scalared signed [4:0] nw9[2:0];
endmodule
